

`timescale 1ns / 100ps

module ThermometerEncoder2 (     

   input  [199:0] thermob,
   output [7:0]   bin

   );

integer k;
reg [199:0] thermo;
reg [7:0]   bin;

always @(thermob) begin

   for (k = 0; k <= 197; k = k + 1)
      thermo[k] <= thermob[k] || thermob[k+1] || thermob[k+2];
	  
   thermo[198] <= thermob[198] || thermob[199];
   thermo[199] <= thermob[199];
   
end

always @(thermo) begin   
    case(thermo)
	  
	  {200'b0     } : bin = 0;
	  {199'b0, 1'b1} : bin = 1;
	  {198'b0, 2'b1} : bin = 2;
	  {197'b0, 3'b1} : bin = 3;  
      {196'b0, 4'b1} : bin = 4;
      {195'b0, 5'b1} : bin = 5;
      {194'b0, 6'b1} : bin = 6;
      {193'b0, 7'b1} : bin = 7;
      {192'b0, 8'b1} : bin = 8;
      {191'b0, 9'b1} : bin = 9;
	  {190'b0, 10'b1} : bin = 10;
	  {189'b0, 11'b1} : bin = 11;
	  {188'b0, 12'b1} : bin = 12;
	  {187'b0, 13'b1} : bin = 13;
	  {186'b0, 14'b1} : bin = 14;
	  {185'b0, 15'b1} : bin = 15;
	  {184'b0, 16'b1} : bin = 16;
	  {183'b0, 17'b1} : bin = 17;
	  {182'b0, 18'b1} : bin = 18;
	  {181'b0, 19'b1} : bin = 19;
	  {180'b0, 20'b1} : bin = 20;
	  {179'b0, 21'b1} : bin = 21;
      {178'b0, 22'b1} : bin = 22;
	  {177'b0, 23'b1} : bin = 23;
	  {176'b0, 24'b1} : bin = 24;
	  {175'b0, 25'b1} : bin = 25;
	  {174'b0, 26'b1} : bin = 26;
	  {173'b0, 27'b1} : bin = 27;
	  {172'b0, 28'b1} : bin = 28;
	  {171'b0, 29'b1} : bin = 29;
	  {170'b0, 30'b1} : bin = 30;
	  {169'b0, 31'b1} : bin = 31;
	  {168'b0, 32'b1} : bin = 32;
	  {167'b0, 33'b1} : bin = 33;
	  {166'b0, 34'b1} : bin = 34;
	  {165'b0, 35'b1} : bin = 35;
	  {164'b0, 36'b1} : bin = 36;
	  {163'b0, 37'b1} : bin = 37;
	  {162'b0, 38'b1} : bin = 38;
	  {161'b0, 39'b1} : bin = 39;
	  {160'b0, 40'b1} : bin = 40;
	  {159'b0, 41'b1} : bin = 41;
	  {158'b0, 42'b1} : bin = 42;
	  {157'b0, 43'b1} : bin = 43;
	  {156'b0, 44'b1} : bin = 44;
      {155'b0, 45'b1} : bin = 45;
	  {154'b0, 46'b1} : bin = 46;
	  {153'b0, 47'b1} : bin = 47;
	  {152'b0, 48'b1} : bin = 48;
	  {151'b0, 49'b1} : bin = 49;
	  {150'b0, 50'b1} : bin = 50;
	  {149'b0, 51'b1} : bin = 51;
	  {148'b0, 52'b1} : bin = 52;
	  {147'b0, 53'b1} : bin = 53;
	  {146'b0, 54'b1} : bin = 54;
	  {145'b0, 55'b1} : bin = 55;
	  {144'b0, 56'b1} : bin = 56;
	  {143'b0, 57'b1} : bin = 57;
	  {142'b0, 58'b1} : bin = 58;
	  {141'b0, 59'b1} : bin = 59;
	  {140'b0, 60'b1} : bin = 60;
	  {139'b0, 61'b1} : bin = 61;
	  {138'b0, 62'b1} : bin = 62;
	  {137'b0, 63'b1} : bin = 63;
	  {136'b0, 64'b1} : bin = 64;
	  {135'b0, 65'b1} : bin = 65;
	  {134'b0, 66'b1} : bin = 66;
	  {133'b0, 67'b1} : bin = 67;
	  {132'b0, 68'b1} : bin = 68;
	  {131'b0, 69'b1} : bin = 69;
	  {130'b0, 70'b1} : bin = 70;
	  {129'b0, 71'b1} : bin = 71;
	  {128'b0, 72'b1} : bin = 72;
	  {127'b0, 73'b1} : bin = 73;
	  {126'b0, 74'b1} : bin = 74;
	  {125'b0, 75'b1} : bin = 75;
	  {124'b0, 76'b1} : bin = 76;
	  {123'b0, 77'b1} : bin = 77;
	  {122'b0, 78'b1} : bin = 78;
	  {121'b0, 79'b1} : bin = 79;
	  {120'b0, 80'b1} : bin = 80;
	  {119'b0, 81'b1} : bin = 81;
	  {118'b0, 82'b1} : bin = 82;
	  {117'b0, 83'b1} : bin = 83;
	  {116'b0, 84'b1} : bin = 84;
	  {115'b0, 85'b1} : bin = 85;
	  {114'b0, 86'b1} : bin = 86;
	  {113'b0, 87'b1} : bin = 87;
	  {112'b0, 88'b1} : bin = 88;
	  {111'b0, 89'b1} : bin = 89;
	  {110'b0, 90'b1} : bin = 90;
	  {109'b0, 91'b1} : bin = 91;
	  {108'b0, 92'b1} : bin = 92;
	  {107'b0, 93'b1} : bin = 93;
	  {106'b0, 94'b1} : bin = 94;
	  {105'b0, 95'b1} : bin = 95;
	  {104'b0, 96'b1} : bin = 96;
	  {103'b0, 97'b1} : bin = 97;
	  {102'b0, 98'b1} : bin = 98;
	  {101'b0, 99'b1} : bin = 99;
	  {100'b0, 100'b1} : bin = 100;
	  {99'b0, 101'b1} : bin = 101;
	  {98'b0, 102'b1} : bin = 102;
	  {97'b0, 103'b1} : bin = 103;
	  {96'b0, 104'b1} : bin = 104;
	  {95'b0, 105'b1} : bin = 105;
	  {94'b0, 106'b1} : bin = 106;
	  {93'b0, 107'b1} : bin = 107;
	  {92'b0, 108'b1} : bin = 108;
	  {91'b0, 109'b1} : bin = 109;
	  {90'b0, 110'b1} : bin = 110;
	  {89'b0, 111'b1} : bin = 111;
	  {88'b0, 112'b1} : bin = 112;
	  {87'b0, 113'b1} : bin = 113;
	  {86'b0, 114'b1} : bin = 114;
	  {85'b0, 115'b1} : bin = 115;
	  {84'b0, 116'b1} : bin = 116;
	  {83'b0, 117'b1} : bin = 117;
	  {82'b0, 118'b1} : bin = 118;
	  {81'b0, 119'b1} : bin = 119;
	  {80'b0, 120'b1} : bin = 120;
	  {79'b0, 121'b1} : bin = 121;
	  {78'b0, 122'b1} : bin = 122;
	  {77'b0, 123'b1} : bin = 123;
	  {76'b0, 124'b1} : bin = 124;
	  {75'b0, 125'b1} : bin = 125;
	  {74'b0, 126'b1} : bin = 126;
	  {73'b0, 127'b1} : bin = 127;
	  {72'b0, 128'b1} : bin = 128;
	  {71'b0, 129'b1} : bin = 129;
	  {70'b0, 130'b1} : bin = 130;
	  {69'b0, 131'b1} : bin = 131;
	  {68'b0, 132'b1} : bin = 132;
	  {67'b0, 133'b1} : bin = 133;
	  {66'b0, 134'b1} : bin = 134;
	  {65'b0, 135'b1} : bin = 135;
	  {64'b0, 136'b1} : bin = 136;
	  {63'b0, 137'b1} : bin = 137;
	  {62'b0, 138'b1} : bin = 138;
	  {61'b0, 139'b1} : bin = 139;
	  {60'b0, 140'b1} : bin = 140;
	  {59'b0, 141'b1} : bin = 141;
	  {58'b0, 142'b1} : bin = 142;
	  {57'b0, 143'b1} : bin = 143;
	  {56'b0, 144'b1} : bin = 144;
	  {55'b0, 145'b1} : bin = 145;
	  {54'b0, 146'b1} : bin = 146;
	  {53'b0, 147'b1} : bin = 147;
	  {52'b0, 148'b1} : bin = 148;
	  {51'b0, 149'b1} : bin = 149;
	  {50'b0, 150'b1} : bin = 150;
	  {49'b0, 151'b1} : bin = 151;
	  {48'b0, 152'b1} : bin = 152;
	  {47'b0, 153'b1} : bin = 153;
	  {46'b0, 154'b1} : bin = 154;
	  {45'b0, 155'b1} : bin = 155;
	  {44'b0, 156'b1} : bin = 156;
	  {43'b0, 157'b1} : bin = 157;
	  {42'b0, 158'b1} : bin = 158;
	  {41'b0, 159'b1} : bin = 159;
	  {40'b0, 160'b1} : bin = 160;
	  {39'b0, 161'b1} : bin = 161;
	  {38'b0, 162'b1} : bin = 162;
	  {37'b0, 163'b1} : bin = 163;
	  {36'b0, 164'b1} : bin = 164;
	  {35'b0, 165'b1} : bin = 165;
	  {34'b0, 166'b1} : bin = 166;
	  {33'b0, 167'b1} : bin = 168;
	  {32'b0, 168'b1} : bin = 169;
	  {31'b0, 169'b1} : bin = 170;
	  {30'b0, 170'b1} : bin = 171;
	  {29'b0, 171'b1} : bin = 172;
	  {28'b0, 172'b1} : bin = 173;
	  {27'b0, 173'b1} : bin = 174;
	  {26'b0, 174'b1} : bin = 175;
	  {25'b0, 175'b1} : bin = 176;
	  {24'b0, 176'b1} : bin = 177;
	  {23'b0, 177'b1} : bin = 178;
	  {22'b0, 178'b1} : bin = 179;
	  {21'b0, 179'b1} : bin = 180;
	  {20'b0, 180'b1} : bin = 181;
	  {19'b0, 181'b1} : bin = 182;
	  {18'b0, 182'b1} : bin = 183;
	  {17'b0, 183'b1} : bin = 184;
	  {16'b0, 184'b1} : bin = 185;
	  {15'b0, 185'b1} : bin = 186;
	  {14'b0, 186'b1} : bin = 187;
	  {13'b0, 187'b1} : bin = 188;
	  {12'b0, 188'b1} : bin = 189;
	  {11'b0, 189'b1} : bin = 190;
	  {10'b0, 190'b1} : bin = 191;
	  {9'b0,  191'b1} : bin = 192;
	  {8'b0,  192'b1} : bin = 193;
	  {7'b0,  193'b1} : bin = 194;
	  {6'b0,  194'b1} : bin = 195;
	  {5'b0,  195'b1} : bin = 196;
	  {4'b0,  196'b1} : bin = 197;
	  {3'b0,  197'b1} : bin = 198;
	  {2'b0,  198'b1} : bin = 199;
	  {1'b0,  199'b1} : bin = 200;
	  {       200'b1} : bin = 200;
	  	  
    endcase
end //always

endmodule
  